* SPICE NETLIST
***************************************

.SUBCKT probe TERM1
.ENDS
***************************************
.SUBCKT thru TERM1 TERM2
.ENDS
***************************************
.SUBCKT v12 TERM1
.ENDS
***************************************
.SUBCKT v20 TERM1
.ENDS
***************************************
.SUBCKT v40 TERM1
.ENDS
***************************************
.SUBCKT ext TERM1
.ENDS
***************************************
.SUBCKT anmvhb G SD B
.ENDS
***************************************
.SUBCKT enmesq G D S B NW
.ENDS
***************************************
.SUBCKT schd PLUS MINUS SUBSTRATE
.ENDS
***************************************
.SUBCKT LDD G S D B
.ENDS
***************************************
.SUBCKT LDDN G S D B
.ENDS
***************************************
.SUBCKT LDDP G S D B
.ENDS
***************************************
.SUBCKT pad74
** N=3 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT my_cap_100p PLUS MINUS
** N=2 EP=2 IP=0 FDC=1
C0 PLUS MINUS L=0.0003 W=0.0003 area=9e-08 peri=0.0012 $[pipc] $X=40510 $Y=1560 $D=47
.ENDS
***************************************
.SUBCKT my_cap_7pF PLUS MINUS
** N=3 EP=2 IP=0 FDC=1
C0 PLUS MINUS L=0.0001 W=8.5e-05 area=8.5e-09 peri=0.00037 $[pipc] $X=1400 $Y=28070 $D=47
.ENDS
***************************************
.SUBCKT schd$$170318892 MINUS SUBSTRATE PLUS
** N=3 EP=3 IP=0 FDC=1
X0 PLUS MINUS SUBSTRATE schd $X=2550 $Y=2550 $D=54
.ENDS
***************************************
.SUBCKT hipor$$168460332 MINUS PLUS
** N=3 EP=2 IP=0 FDC=1
R0 MINUS PLUS L=4e-06 W=4e-06 nsq=1 $[hipor] $X=0 $Y=0 $D=41
.ENDS
***************************************
.SUBCKT dickson_schd_N_caplay gnd! rf_mod mod_gate vdd rf_detect rf_in
** N=35 EP=6 IP=120 FDC=40
C0 rf_detect gnd! L=0.0001 W=8.5e-05 area=8.5e-09 peri=0.00037 $[pipc] $X=472140 $Y=217100 $D=47
M1 rf_mod mod_gate gnd! gnd! nenm L=6e-07 W=5e-06 $X=180120 $Y=286320 $D=77
X9 vdd gnd! my_cap_100p $T=584130 215550 0 0 $X=584130 $Y=215708
X10 28 rf_in my_cap_7pF $T=209680 422880 0 0 $X=209680 $Y=439380
X11 29 gnd! my_cap_7pF $T=227820 330170 1 0 $X=227820 $Y=215700
X12 30 rf_in my_cap_7pF $T=326330 422880 0 0 $X=326330 $Y=439380
X13 31 gnd! my_cap_7pF $T=349570 330170 1 0 $X=349570 $Y=215700
X14 32 rf_in my_cap_7pF $T=447280 422880 0 0 $X=447280 $Y=439380
X15 28 gnd! gnd! schd$$170318892 $T=254100 369260 1 180 $X=240600 $Y=369260
X16 29 gnd! 28 schd$$170318892 $T=278950 402210 0 180 $X=265450 $Y=369210
X17 30 gnd! 29 schd$$170318892 $T=302760 369260 1 180 $X=289260 $Y=369260
X18 31 gnd! 30 schd$$170318892 $T=327820 402210 0 180 $X=314320 $Y=369210
X19 32 gnd! 31 schd$$170318892 $T=351960 369260 1 180 $X=338460 $Y=369260
X20 rf_detect gnd! 32 schd$$170318892 $T=376960 402210 0 180 $X=363460 $Y=369210
X21 vdd gnd! 32 schd$$170318892 $T=404890 402210 0 180 $X=391390 $Y=369210
X22 mod_gate 6 hipor$$168460332 $T=213410 117010 0 0 $X=212410 $Y=115810
X23 5 3 hipor$$168460332 $T=213410 124610 0 0 $X=212410 $Y=123410
X24 3 8 hipor$$168460332 $T=213410 132210 0 0 $X=212410 $Y=131010
X25 7 4 hipor$$168460332 $T=213410 139810 0 0 $X=212410 $Y=138610
X26 4 9 hipor$$168460332 $T=213410 147410 0 0 $X=212410 $Y=146210
X27 12 6 hipor$$168460332 $T=221010 117010 0 0 $X=220010 $Y=115810
X28 5 15 hipor$$168460332 $T=221010 124610 0 0 $X=220010 $Y=123410
X29 11 8 hipor$$168460332 $T=221010 132210 0 0 $X=220010 $Y=131010
X30 7 13 hipor$$168460332 $T=221010 139810 0 0 $X=220010 $Y=138610
X31 14 9 hipor$$168460332 $T=221010 147410 0 0 $X=220010 $Y=146210
X32 12 17 hipor$$168460332 $T=228610 117010 0 0 $X=227610 $Y=115810
X33 18 15 hipor$$168460332 $T=228610 124610 0 0 $X=227610 $Y=123410
X34 11 19 hipor$$168460332 $T=228610 132210 0 0 $X=227610 $Y=131010
X35 20 13 hipor$$168460332 $T=228610 139810 0 0 $X=227610 $Y=138610
X36 14 16 hipor$$168460332 $T=228610 147410 0 0 $X=227610 $Y=146210
X37 24 17 hipor$$168460332 $T=236210 117010 0 0 $X=235210 $Y=115810
X38 18 21 hipor$$168460332 $T=236210 124610 0 0 $X=235210 $Y=123410
X39 23 19 hipor$$168460332 $T=236210 132210 0 0 $X=235210 $Y=131010
X40 20 22 hipor$$168460332 $T=236210 139810 0 0 $X=235210 $Y=138610
X41 25 16 hipor$$168460332 $T=236210 147410 0 0 $X=235210 $Y=146210
X42 24 26 hipor$$168460332 $T=243810 117010 0 0 $X=242810 $Y=115810
X43 26 21 hipor$$168460332 $T=243810 124610 0 0 $X=242810 $Y=123410
X44 23 27 hipor$$168460332 $T=243810 132210 0 0 $X=242810 $Y=131010
X45 27 22 hipor$$168460332 $T=243810 139810 0 0 $X=242810 $Y=138610
X46 25 gnd! hipor$$168460332 $T=243810 147410 0 0 $X=242810 $Y=146210
.ENDS
***************************************
